-- Company: Taksun
-- Engineer: Hosseinali 
-- Description: This design is written with the help of https://github.com/iamhosseinali/SINE_WAVE_VHDL_GENERATOR repo
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity Sine_Wave_Gen is
generic (
    IP_INPUT_FREQUENCY                  : integer := 100000000; --- in Hz
    DEFAULT_OUTPUT_SIGNAL_FREQUENCY     : integer := 50        --- in Hz, max = M_AXIS_ACLK/2048.
);
Port (
    M_AXIS_ACLK    : in STD_LOGIC;
    M_AXIS_ARESETN : in STD_LOGIC; 
    M_AXIS_tDATA   : out std_logic_vector(7 downto 0);
    M_AXIS_tVALID  : out std_logic;
    Config         : in std_logic_vector(31 downto 0) -- (31) valid_flag, (30:0) IP_INPUT_FREQUENCY/OUTPUT_SIGNAL_FREQUENCY/1024;
);
end Sine_Wave_Gen;

architecture Behavioral of Sine_Wave_Gen is

constant SIN_TABLE_Length          : integer := 1024;
constant SIN_DATA_WIDTH            : integer := 8;
type SIN_TABLEType is array(0 to SIN_TABLE_Length-1) of integer;
constant SIN_TABLE : SIN_TABLEType :=(0,0,1,2,3,3,4,5,6,7,7,8,9,10,10,11,12,13,14,14,15,16,17,18,18,19,20,21,21,22,23,24,24,25,26,27,28,28,29,30,31,31,32,33,34,34,35,36,37,37,38,39,40,40,41,42,43,43,44,45,46,46,47,48,48,49,50,51,51,52,53,54,54,55,56,56,57,58,58,59,60,61,61,62,63,63,64,65,65,66,67,67,68,69,69,70,71,71,72,73,73,74,74,75,76,76,77,78,78,79,79,80,81,81,82,83,83,84,84,85,85,86,87,87,88,88,89,89,90,91,91,92,92,93,93,94,94,95,95,96,96,97,97,98,98,99,99,100,100,101,101,102,102,103,103,104,104,105,105,105,106,106,107,107,108,108,108,109,109,110,110,110,111,111,112,112,112,113,113,113,114,114,115,115,115,116,116,116,117,117,117,117,118,118,118,119,119,119,119,120,120,120,121,121,121,121,122,122,122,122,122,123,123,123,123,123,124,124,124,124,124,125,125,125,125,125,125,125,126,126,126,126,126,126,126,126,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,127,126,126,126,126,126,126,126,126,125,125,125,125,125,125,125,124,124,124,124,124,123,123,123,123,123,122,122,122,122,122,121,121,121,121,120,120,120,119,119,119,119,118,118,118,117,117,117,117,116,116,116,115,115,115,114,114,113,113,113,112,112,112,111,111,110,110,110,109,109,108,108,108,107,107,106,106,105,105,105,104,104,103,103,102,102,101,101,100,100,99,99,98,98,97,97,96,96,95,95,94,94,93,93,92,92,91,91,90,89,89,88,88,87,87,86,85,85,84,84,83,83,82,81,81,80,79,79,78,78,77,76,76,75,74,74,73,73,72,71,71,70,69,69,68,67,67,66,65,65,64,63,63,62,61,61,60,59,58,58,57,56,56,55,54,54,53,52,51,51,50,49,48,48,47,46,46,45,44,43,43,42,41,40,40,39,38,37,37,36,35,34,34,33,32,31,31,30,29,28,28,27,26,25,24,24,23,22,21,21,20,19,18,18,17,16,15,14,14,13,12,11,10,10,9,8,7,7,6,5,4,3,3,2,1,0,0,0,-1,-2,-3,-3,-4,-5,-6,-7,-7,-8,-9,-10,-10,-11,-12,-13,-14,-14,-15,-16,-17,-18,-18,-19,-20,-21,-21,-22,-23,-24,-24,-25,-26,-27,-28,-28,-29,-30,-31,-31,-32,-33,-34,-34,-35,-36,-37,-37,-38,-39,-40,-40,-41,-42,-43,-43,-44,-45,-46,-46,-47,-48,-48,-49,-50,-51,-51,-52,-53,-54,-54,-55,-56,-56,-57,-58,-58,-59,-60,-61,-61,-62,-63,-63,-64,-65,-65,-66,-67,-67,-68,-69,-69,-70,-71,-71,-72,-73,-73,-74,-74,-75,-76,-76,-77,-78,-78,-79,-79,-80,-81,-81,-82,-83,-83,-84,-84,-85,-85,-86,-87,-87,-88,-88,-89,-89,-90,-91,-91,-92,-92,-93,-93,-94,-94,-95,-95,-96,-96,-97,-97,-98,-98,-99,-99,-100,-100,-101,-101,-102,-102,-103,-103,-104,-104,-105,-105,-105,-106,-106,-107,-107,-108,-108,-108,-109,-109,-110,-110,-110,-111,-111,-112,-112,-112,-113,-113,-113,-114,-114,-115,-115,-115,-116,-116,-116,-117,-117,-117,-117,-118,-118,-118,-119,-119,-119,-119,-120,-120,-120,-121,-121,-121,-121,-122,-122,-122,-122,-122,-123,-123,-123,-123,-123,-124,-124,-124,-124,-124,-125,-125,-125,-125,-125,-125,-125,-126,-126,-126,-126,-126,-126,-126,-126,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-127,-126,-126,-126,-126,-126,-126,-126,-126,-125,-125,-125,-125,-125,-125,-125,-124,-124,-124,-124,-124,-123,-123,-123,-123,-123,-122,-122,-122,-122,-122,-121,-121,-121,-121,-120,-120,-120,-119,-119,-119,-119,-118,-118,-118,-117,-117,-117,-117,-116,-116,-116,-115,-115,-115,-114,-114,-113,-113,-113,-112,-112,-112,-111,-111,-110,-110,-110,-109,-109,-108,-108,-108,-107,-107,-106,-106,-105,-105,-105,-104,-104,-103,-103,-102,-102,-101,-101,-100,-100,-99,-99,-98,-98,-97,-97,-96,-96,-95,-95,-94,-94,-93,-93,-92,-92,-91,-91,-90,-89,-89,-88,-88,-87,-87,-86,-85,-85,-84,-84,-83,-83,-82,-81,-81,-80,-79,-79,-78,-78,-77,-76,-76,-75,-74,-74,-73,-73,-72,-71,-71,-70,-69,-69,-68,-67,-67,-66,-65,-65,-64,-63,-63,-62,-61,-61,-60,-59,-58,-58,-57,-56,-56,-55,-54,-54,-53,-52,-51,-51,-50,-49,-48,-48,-47,-46,-46,-45,-44,-43,-43,-42,-41,-40,-40,-39,-38,-37,-37,-36,-35,-34,-34,-33,-32,-31,-31,-30,-29,-28,-28,-27,-26,-25,-24,-24,-23,-22,-21,-21,-20,-19,-18,-18,-17,-16,-15,-14,-14,-13,-12,-11,-10,-10,-9,-8,-7,-7,-6,-5,-4,-3,-3,-2,-1,0);
attribute ram_style : string;
attribute ram_style of SIN_TABLE : constant is "block";
constant def_indx_cycle            : integer := IP_INPUT_FREQUENCY/DEFAULT_OUTPUT_SIGNAL_FREQUENCY/SIN_TABLE_Length;
signal indx_cycle                  : unsigned(30 downto 0) := to_unsigned(def_indx_cycle,31);
signal sin_indx                    : unsigned(9 downto 0) := (others=>'0');
signal cnt                         : unsigned(31 downto 0) := (others=>'0');
signal valid_flag_int              : std_logic := '0';  
signal Config_int                  : std_logic_vector(31 downto 0) := (others=>'0');

begin

process(M_AXIS_ACLK)
begin
    if rising_edge(M_AXIS_ACLK) then
       if (M_AXIS_ARESETN='0') then
           cnt             <= (others=>'0');
           sin_indx        <= (others=>'0');
           M_AXIS_tVALID   <= '0';
           indx_cycle      <= to_unsigned(def_indx_cycle,31);
       else
            Config_int         <= Config;
            cnt                <= cnt+1;
            indx_cycle  <= to_unsigned(def_indx_cycle,31);
            if(Config(31) = '1') then
                indx_cycle  <= unsigned(Config_int(30 downto 0)); 
            end if;
            M_AXIS_tVALID   <= '0';
            if(cnt=indx_cycle)then
                cnt        <= (others=>'0');
                sin_indx   <= sin_indx+1;
                if(sin_indx=SIN_TABLE_Length-1) then
                    sin_indx       <= (others=>'0');
                end if;
                M_AXIS_tVALID  <= '1';
                M_AXIS_tDATA   <= std_logic_vector(to_signed(SIN_TABLE(to_integer(sin_indx)),SIN_DATA_WIDTH));
            end if;
            if((Config_int(31) = '0' and Config(31) = '1') or (Config_int(31) = '1' and Config(31) = '0')) then 
                cnt        <= (others=>'0');
            end if;
       end if;
    end if;
end process;
end Behavioral;
